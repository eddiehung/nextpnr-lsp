module blinky (
    input  clki,
    output led1,
);
    assign led1 = clki;
endmodule
